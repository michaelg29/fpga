class test_class;

static function void print_hello();
    $display("Hello, world!\n");
endfunction

endclass