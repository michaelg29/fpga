package test_pkg;

    // import uvm_pkg::*;

    // `include "uvm_macros.svh";
    `include "test_class.svh";

endpackage