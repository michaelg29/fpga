package test_pkg;

    //import uvm_pkg::*;

    `include "test_class.svh";

endpackage